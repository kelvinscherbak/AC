CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
40 97 1560 833
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
40 97 1560 833
177209362 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 560 107 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 520 108 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 295 335 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 296 290 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6153 0 0
0
0
9 Inverter~
13 590 238 0 2 22
0 7 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 7 0
1 U
5394 0 0
0
0
9 Inverter~
13 590 295 0 2 22
0 8 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 7 0
1 U
7734 0 0
0
0
9 Inverter~
13 578 323 0 2 22
0 8 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 7 0
1 U
9914 0 0
0
0
9 Inverter~
13 589 336 0 2 22
0 7 12
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
3747 0 0
0
0
14 Logic Display~
6 898 239 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
9 2-In AND~
219 411 320 0 3 22
0 3 2 4
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7931 0 0
0
0
8 2-In OR~
219 405 267 0 3 22
0 3 2 5
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9325 0 0
0
0
9 2-In XOR~
219 406 209 0 3 22
0 3 2 6
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
8903 0 0
0
0
14 Logic Display~
6 450 110 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
9 2-In AND~
219 380 146 0 3 22
0 3 2 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3363 0 0
0
0
8 4-In OR~
219 822 270 0 5 22
0 17 16 15 14 13
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 1996002869
65 0 0 0 2 1 3 0
1 U
7668 0 0
0
0
9 3-In AND~
219 645 337 0 4 22
0 11 12 4 14
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
4718 0 0
0
0
9 3-In AND~
219 646 295 0 4 22
0 7 9 5 15
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 1 0
1 U
3874 0 0
0
0
9 3-In AND~
219 648 248 0 4 22
0 10 8 6 16
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 1 0
1 U
6671 0 0
0
0
9 3-In AND~
219 648 200 0 4 22
0 7 8 6 17
0
0 0 624 0
6 74LS11
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 1 0
1 U
3789 0 0
0
0
30
2 0 2 0 0 4096 0 12 0 0 29 2
390 218
355 218
1 0 3 0 0 4096 0 12 0 0 28 2
390 200
324 200
3 3 4 0 0 12416 0 10 16 0 0 4
432 320
471 320
471 346
621 346
3 3 5 0 0 4224 0 17 11 0 0 4
622 304
471 304
471 267
438 267
3 0 6 0 0 4224 0 18 0 0 6 3
624 257
483 257
483 229
3 3 6 0 0 0 0 12 19 0 0 6
439 209
483 209
483 229
483 229
483 209
624 209
1 0 7 0 0 4096 0 19 0 0 18 2
624 191
520 191
2 0 8 0 0 4096 0 19 0 0 15 2
624 200
563 200
1 0 7 0 0 0 0 17 0 0 18 2
622 286
520 286
2 2 9 0 0 4224 0 17 6 0 0 2
622 295
611 295
2 1 10 0 0 8320 0 5 18 0 0 3
611 238
611 239
624 239
2 0 8 0 0 0 0 18 0 0 15 2
624 248
563 248
1 0 7 0 0 0 0 5 0 0 18 2
575 238
520 238
1 0 8 0 0 0 0 6 0 0 15 2
575 295
563 295
1 1 8 0 0 8320 0 1 7 0 0 3
560 119
563 119
563 323
2 1 11 0 0 12416 0 7 16 0 0 4
599 323
606 323
606 328
621 328
2 2 12 0 0 8320 0 8 16 0 0 3
610 336
610 337
621 337
1 1 7 0 0 4224 0 2 8 0 0 3
520 120
520 336
574 336
1 5 13 0 0 8320 0 9 15 0 0 3
898 257
898 270
855 270
4 4 14 0 0 12416 0 15 16 0 0 4
805 284
764 284
764 337
666 337
3 4 15 0 0 4224 0 15 17 0 0 4
805 275
712 275
712 295
667 295
4 2 16 0 0 4224 0 18 15 0 0 4
669 248
739 248
739 266
805 266
1 4 17 0 0 12416 0 15 19 0 0 4
805 257
783 257
783 200
669 200
1 0 3 0 0 4096 0 11 0 0 28 2
392 258
324 258
2 0 2 0 0 4096 0 11 0 0 29 2
392 276
355 276
1 0 3 0 0 0 0 10 0 0 28 3
387 311
324 311
324 287
2 0 2 0 0 0 0 10 0 0 29 2
387 329
355 329
1 1 3 0 0 8320 0 14 4 0 0 4
356 137
324 137
324 290
308 290
2 1 2 0 0 8320 0 14 3 0 0 4
356 155
355 155
355 335
307 335
1 3 18 0 0 8320 0 13 14 0 0 3
450 128
450 146
401 146
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
430 59 478 83
438 67 478 83
5 c.out
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
872 188 912 212
882 196 914 212
4 C.in
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
